`define CLK_PERIOD_NS  40  // 25 MHz
`define DEBOUNCE_MASK_PERIOD_MS 20 

